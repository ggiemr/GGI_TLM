Ngspice template file for GGI_TLM - ngspice linked simulation
*
* GGI_TLM link port    1 using nodes    1 and   0
*
* Voltage source with series resistance: equivalent circuit of TLM link
 Vtlm1        1001           0  DC  0.0
 Rtlm1        1001           1  #Z0_TLM
* 
* Model to be included in the GGI_TLM simulation
* GGI_TLM link port    2 using nodes    2 and   3
*
* Voltage source with series resistance: equivalent circuit of TLM link
 Vtlm2        1002           3  DC  0.0
 Rtlm2        1002           2  #Z0_TLM
* 
* Model to be included in the GGI_TLM simulation
* GGI_TLM link port    3 using nodes    3 and   0
*
* Voltage source with series resistance: equivalent circuit of TLM link
 Vtlm3        1003           0  DC  0.0
 Rtlm3        1003           3  #Z0_TLM
* 
* Model to be included in the GGI_TLM simulation

* Model to be included in the GGI_TLM simulation for port 1, connected to node 1
* in this case a voltage source with series resistance
Rs1     2001   1   1000.0
Vs1     2001   0   EXP( 0.0     1.0    0.000000E+00    1.000000E-010    1.200000E-08    1.000000E-010 )
*
* Model to be included in the GGI_TLM simulation for port 1, connected to nodes 2 and 3
* in this case a diode with series resistance
Rl23      2   3   1000.0
* Model to be included in the GGI_TLM simulation for port 2, connected to node 3 and 0
* in this case a diode with series resistance
Rl30      3   0   1000.0
*
Rl20      2   0   2000.0
*

*
* Control for transient simulation
.TRAN #dt_ngspice  #tmax_ngspice  #dt_ngspice  UIC
*
.END
