test circuit file for circuit elements to be embedded in GGI_TLM
*
* The test circuit is in two parts, the source end model and the load end model.
* The source end model consists of a pulse voltage source in series with a 100 ohm resistance: GGI_TLM interface connected to node 1.
* The load end model consists of a diode in series with a 100 ohm resistance: GGI_TLM interface connected to node 2.
* 1e-12  0.026   1e-10 1e-18 # Diode model parameters in reference TLM solution: Is and nVt values series_resistance junction_capacitance
*
* Voltage source with series resistance: equivalent circuit of TLM link
Vtlm1  1002   0   DC  0.0
Rtlm1  1002   1   #Z0_TLM
* 
* Model to be included in the GGI_TLM simulation in this case a voltage source with series resistance
Rs1     1003   1   100.0
Vs1     1003   0   EXP( 0.0     1.0    0.000000E+00    2.000000E-09    1.200000E-08    2.000000E-09 )
*
* Voltage source with series resistance: equivalent circuit of TLM link
Vtlm2  1022   0   DC  0.0
Rtlm2  1022   2   #Z0_TLM
* 
* Model to be included in the GGI_TLM simulation
Diode2   1023   2   Dmod
Rl2     1023   0   100.0
.model DMOD D ( is=1e-12 )
*
Vbreak time_node 0 DC 0.0
*
* Control for transient simulation
.tran #dt_ngspice  #tmax_ngspice  #dt_ngspice
*
.end
