Ngspice template file for GGI_TLM - ngspice linked simulation
*
* GGI_TLM link through node      1
*
* Voltage source with series resistance: equivalent circuit of TLM link
 Vtlm1        1001           0  DC  0.0
 Rtlm1        1001           1  #Z0_TLM
* 
* Model to be included in the GGI_TLM simulation
* GGI_TLM link through node      2
*
* Voltage source with series resistance: equivalent circuit of TLM link
 Vtlm2        1002           0  DC  0.0
 Rtlm2        1002           2  #Z0_TLM
* 
* Model to be included in the GGI_TLM simulation

* Model to be included in the GGI_TLM simulation for port 1, connected to node 1
* in this case a voltage source with series resistance
Rs1     2001   1   100.0
Vs1     2001   0   EXP( 0.0     1.0    0.000000E+00    2.000000E-010    1.200000E-09    2.000000E-010 )
*
* Model to be included in the GGI_TLM simulation for port 2, connected to node 2
* in this case a diode with series resistance
Diode2   2002   2   Dmod
Rl2      2002   0   100.0
.model DMOD D ( is=1e-12 )
*

*
* Control for transient simulation
.TRAN #dt_ngspice  #tmax_ngspice  #dt_ngspice  UIC
*
.END
