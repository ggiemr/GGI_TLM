test circuit file for circuit elements to be embedded in GGI_TLM
* The test circuit consists of a diode model
* 1e-12  0.026   1e-10 1e-18 # Diode model parameters in reference TLM solution: Is and nVt values series_resistance junction_capacitance
*
* Load end model: ngspice handles the diode in series with 100 ohm resistance
* The voltage transferred in V(1)
*
* Voltage source with series resistance: equivalent circuit of TLM link
Vtlm2  1002   0   DC  0.0
Rtlm2  1002   1   #Z0_TLM
* 
* Model of impedance to be included in the GGI_TLM simulation
Diode  1003   1   Dmod
Rl     1003   0   100.0
*
.model DMOD D ( is=1e-12 )
*
* Control for transient simulation
.tran #dt_ngspice  #tmax_ngspice  #dt_ngspice
*
.end
